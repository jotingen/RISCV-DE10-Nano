package LC3_pkg;

typedef enum {
  IFU_FETCH,
  IDU_DECODE,
  ALU_EXECUTE
} state;

endpackage
