package riscv_pkg;


endpackage
