
module soc_system (
	clk_clk,
	ddr3_clk_clk);	

	input		clk_clk;
	output		ddr3_clk_clk;
endmodule
