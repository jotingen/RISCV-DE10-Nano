// soc_system.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module soc_system (
		input  wire  clk_clk,      //      clk.clk
		output wire  ddr3_clk_clk  // ddr3_clk.clk
	);

	soc_system_ddr3 ddr3 (
	);

	soc_system_pll pll (
		.refclk   (clk_clk),      //  refclk.clk
		.rst      (),             //   reset.reset
		.outclk_0 (ddr3_clk_clk), // outclk0.clk
		.locked   ()              // (terminated)
	);

endmodule
